
-- Company: 			Dossytronics
-- Engineer: 			Dominic Beesley
-- 
-- Create Date:    		9/3/2018
-- Design Name: 
-- Module Name:    		work.board_config_pack
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 		shared types
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------

library ieee;
use IEEE.math_real.all;

package sim_SYS_pack is
	type sim_SYS_type is (SIM_SYS_BBC, SIM_SYS_ELK);



end sim_SYS_pack;


package body sim_SYS_pack is

end sim_SYS_pack;
