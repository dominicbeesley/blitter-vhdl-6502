library ieee;
use IEEE.math_real.all;

package fb_CPU_pack is
	type cpu_type is (CPU_6x09, CPU_6502, CPU_65C02, CPU_65816, CPU_Z80, CPU_68008);

end fb_CPU_pack;


package body fb_CPU_pack is

end fb_CPU_pack;
