library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity saa5050_rom_dual_port is
    generic (
        ADDR_WIDTH       : integer := 12;
        DATA_WIDTH       : integer := 8
    );
    port(
        clock    : in  std_logic;
        addressA : in  std_logic_vector(11 downto 0);
        QA       : out std_logic_vector(7 downto 0);
        addressB : in  std_logic_vector(11 downto 0);
        QB       : out std_logic_vector(7 downto 0)
  );
end saa5050_rom_dual_port;

architecture RTL of saa5050_rom_dual_port is

signal	r_switch : std_logic := '0';

begin

p:process(CLOCK)
variable A:std_logic_vector(11 downto 0);
variable Q:std_logic_vector(5 downto 0);
variable TOP:std_logic;
begin

	if (rising_edge(CLOCK)) then
		if (r_switch = '0') then
			A := addressA;
		else
			A := addressB;
		end if;

		case ("0" & A(10 downto 0)) is

-- CH=21 "!"
         when x"211" => Q := "000100";
         when x"212" => Q := "000100";
         when x"213" => Q := "000100";
         when x"214" => Q := "000100";
         when x"215" => Q := "000100";
         when x"217" => Q := "000100";


-- CH=22 """
         when x"221" => Q := "001010";
         when x"222" => Q := "001010";
         when x"223" => Q := "001010";


-- CH=23 "#"
         when x"231" => Q := "000110";
         when x"232" => Q := "001001";
         when x"233" => Q := "001000";
         when x"234" => Q := "011100";
         when x"235" => Q := "001000";
         when x"236" => Q := "001000";
         when x"237" => Q := "011111";


-- CH=24 "$"
         when x"241" => Q := "001110";
         when x"242" => Q := "010101";
         when x"243" => Q := "010100";
         when x"244" => Q := "001110";
         when x"245" => Q := "000101";
         when x"246" => Q := "010101";
         when x"247" => Q := "001110";


-- CH=25 "%"
         when x"251" => Q := "011000";
         when x"252" => Q := "011001";
         when x"253" => Q := "000010";
         when x"254" => Q := "000100";
         when x"255" => Q := "001000";
         when x"256" => Q := "010011";
         when x"257" => Q := "000011";


-- CH=26 "&"
         when x"261" => Q := "001000";
         when x"262" => Q := "010100";
         when x"263" => Q := "010100";
         when x"264" => Q := "001000";
         when x"265" => Q := "010101";
         when x"266" => Q := "010010";
         when x"267" => Q := "001101";


-- CH=27 "'"
         when x"271" => Q := "000100";
         when x"272" => Q := "000100";
         when x"273" => Q := "000100";


-- CH=28 "("
         when x"281" => Q := "000010";
         when x"282" => Q := "000100";
         when x"283" => Q := "001000";
         when x"284" => Q := "001000";
         when x"285" => Q := "001000";
         when x"286" => Q := "000100";
         when x"287" => Q := "000010";


-- CH=29 ")"
         when x"291" => Q := "001000";
         when x"292" => Q := "000100";
         when x"293" => Q := "000010";
         when x"294" => Q := "000010";
         when x"295" => Q := "000010";
         when x"296" => Q := "000100";
         when x"297" => Q := "001000";


-- CH=2A "*"
         when x"2A1" => Q := "000100";
         when x"2A2" => Q := "010101";
         when x"2A3" => Q := "001110";
         when x"2A4" => Q := "000100";
         when x"2A5" => Q := "001110";
         when x"2A6" => Q := "010101";
         when x"2A7" => Q := "000100";


-- CH=2B "+"
         when x"2B2" => Q := "000100";
         when x"2B3" => Q := "000100";
         when x"2B4" => Q := "011111";
         when x"2B5" => Q := "000100";
         when x"2B6" => Q := "000100";


-- CH=2C ","
         when x"2C6" => Q := "000100";
         when x"2C7" => Q := "000100";
         when x"2C8" => Q := "001000";


-- CH=2D "-"
         when x"2D4" => Q := "001110";


-- CH=2E "."
         when x"2E7" => Q := "000100";


-- CH=2F "/"
         when x"2F2" => Q := "000001";
         when x"2F3" => Q := "000010";
         when x"2F4" => Q := "000100";
         when x"2F5" => Q := "001000";
         when x"2F6" => Q := "010000";


-- CH=30 "0"
         when x"301" => Q := "000100";
         when x"302" => Q := "001010";
         when x"303" => Q := "010001";
         when x"304" => Q := "010001";
         when x"305" => Q := "010001";
         when x"306" => Q := "001010";
         when x"307" => Q := "000100";


-- CH=31 "1"
         when x"311" => Q := "000100";
         when x"312" => Q := "001100";
         when x"313" => Q := "000100";
         when x"314" => Q := "000100";
         when x"315" => Q := "000100";
         when x"316" => Q := "000100";
         when x"317" => Q := "001110";


-- CH=32 "2"
         when x"321" => Q := "001110";
         when x"322" => Q := "010001";
         when x"323" => Q := "000001";
         when x"324" => Q := "000110";
         when x"325" => Q := "001000";
         when x"326" => Q := "010000";
         when x"327" => Q := "011111";


-- CH=33 "3"
         when x"331" => Q := "011111";
         when x"332" => Q := "000001";
         when x"333" => Q := "000010";
         when x"334" => Q := "000110";
         when x"335" => Q := "000001";
         when x"336" => Q := "010001";
         when x"337" => Q := "001110";


-- CH=34 "4"
         when x"341" => Q := "000010";
         when x"342" => Q := "000110";
         when x"343" => Q := "001010";
         when x"344" => Q := "010010";
         when x"345" => Q := "011111";
         when x"346" => Q := "000010";
         when x"347" => Q := "000010";


-- CH=35 "5"
         when x"351" => Q := "011111";
         when x"352" => Q := "010000";
         when x"353" => Q := "011110";
         when x"354" => Q := "000001";
         when x"355" => Q := "000001";
         when x"356" => Q := "010001";
         when x"357" => Q := "001110";


-- CH=36 "6"
         when x"361" => Q := "000110";
         when x"362" => Q := "001000";
         when x"363" => Q := "010000";
         when x"364" => Q := "011110";
         when x"365" => Q := "010001";
         when x"366" => Q := "010001";
         when x"367" => Q := "001110";


-- CH=37 "7"
         when x"371" => Q := "011111";
         when x"372" => Q := "000001";
         when x"373" => Q := "000010";
         when x"374" => Q := "000100";
         when x"375" => Q := "001000";
         when x"376" => Q := "001000";
         when x"377" => Q := "001000";


-- CH=38 "8"
         when x"381" => Q := "001110";
         when x"382" => Q := "010001";
         when x"383" => Q := "010001";
         when x"384" => Q := "001110";
         when x"385" => Q := "010001";
         when x"386" => Q := "010001";
         when x"387" => Q := "001110";


-- CH=39 "9"
         when x"391" => Q := "001110";
         when x"392" => Q := "010001";
         when x"393" => Q := "010001";
         when x"394" => Q := "001111";
         when x"395" => Q := "000001";
         when x"396" => Q := "000010";
         when x"397" => Q := "001100";


-- CH=3A ":"
         when x"3A3" => Q := "000100";
         when x"3A7" => Q := "000100";


-- CH=3B ";"
         when x"3B3" => Q := "000100";
         when x"3B6" => Q := "000100";
         when x"3B7" => Q := "000100";
         when x"3B8" => Q := "001000";


-- CH=3C "<"
         when x"3C1" => Q := "000010";
         when x"3C2" => Q := "000100";
         when x"3C3" => Q := "001000";
         when x"3C4" => Q := "010000";
         when x"3C5" => Q := "001000";
         when x"3C6" => Q := "000100";
         when x"3C7" => Q := "000010";


-- CH=3D "="
         when x"3D3" => Q := "011111";
         when x"3D5" => Q := "011111";


-- CH=3E ">"
         when x"3E1" => Q := "001000";
         when x"3E2" => Q := "000100";
         when x"3E3" => Q := "000010";
         when x"3E4" => Q := "000001";
         when x"3E5" => Q := "000010";
         when x"3E6" => Q := "000100";
         when x"3E7" => Q := "001000";


-- CH=3F "?"
         when x"3F1" => Q := "001110";
         when x"3F2" => Q := "010001";
         when x"3F3" => Q := "000010";
         when x"3F4" => Q := "000100";
         when x"3F5" => Q := "000100";
         when x"3F7" => Q := "000100";


-- CH=40 "@"
         when x"401" => Q := "001110";
         when x"402" => Q := "010001";
         when x"403" => Q := "010111";
         when x"404" => Q := "010101";
         when x"405" => Q := "010111";
         when x"406" => Q := "010000";
         when x"407" => Q := "001110";


-- CH=41 "A"
         when x"411" => Q := "000100";
         when x"412" => Q := "001010";
         when x"413" => Q := "010001";
         when x"414" => Q := "010001";
         when x"415" => Q := "011111";
         when x"416" => Q := "010001";
         when x"417" => Q := "010001";


-- CH=42 "B"
         when x"421" => Q := "011110";
         when x"422" => Q := "010001";
         when x"423" => Q := "010001";
         when x"424" => Q := "011110";
         when x"425" => Q := "010001";
         when x"426" => Q := "010001";
         when x"427" => Q := "011110";


-- CH=43 "C"
         when x"431" => Q := "001110";
         when x"432" => Q := "010001";
         when x"433" => Q := "010000";
         when x"434" => Q := "010000";
         when x"435" => Q := "010000";
         when x"436" => Q := "010001";
         when x"437" => Q := "001110";


-- CH=44 "D"
         when x"441" => Q := "011110";
         when x"442" => Q := "010001";
         when x"443" => Q := "010001";
         when x"444" => Q := "010001";
         when x"445" => Q := "010001";
         when x"446" => Q := "010001";
         when x"447" => Q := "011110";


-- CH=45 "E"
         when x"451" => Q := "011111";
         when x"452" => Q := "010000";
         when x"453" => Q := "010000";
         when x"454" => Q := "011110";
         when x"455" => Q := "010000";
         when x"456" => Q := "010000";
         when x"457" => Q := "011111";


-- CH=46 "F"
         when x"461" => Q := "011111";
         when x"462" => Q := "010000";
         when x"463" => Q := "010000";
         when x"464" => Q := "011110";
         when x"465" => Q := "010000";
         when x"466" => Q := "010000";
         when x"467" => Q := "010000";


-- CH=47 "G"
         when x"471" => Q := "001110";
         when x"472" => Q := "010001";
         when x"473" => Q := "010000";
         when x"474" => Q := "010000";
         when x"475" => Q := "010011";
         when x"476" => Q := "010001";
         when x"477" => Q := "001111";


-- CH=48 "H"
         when x"481" => Q := "010001";
         when x"482" => Q := "010001";
         when x"483" => Q := "010001";
         when x"484" => Q := "011111";
         when x"485" => Q := "010001";
         when x"486" => Q := "010001";
         when x"487" => Q := "010001";


-- CH=49 "I"
         when x"491" => Q := "001110";
         when x"492" => Q := "000100";
         when x"493" => Q := "000100";
         when x"494" => Q := "000100";
         when x"495" => Q := "000100";
         when x"496" => Q := "000100";
         when x"497" => Q := "001110";


-- CH=4A "J"
         when x"4A1" => Q := "000001";
         when x"4A2" => Q := "000001";
         when x"4A3" => Q := "000001";
         when x"4A4" => Q := "000001";
         when x"4A5" => Q := "000001";
         when x"4A6" => Q := "010001";
         when x"4A7" => Q := "001110";


-- CH=4B "K"
         when x"4B1" => Q := "010001";
         when x"4B2" => Q := "010010";
         when x"4B3" => Q := "010100";
         when x"4B4" => Q := "011000";
         when x"4B5" => Q := "010100";
         when x"4B6" => Q := "010010";
         when x"4B7" => Q := "010001";


-- CH=4C "L"
         when x"4C1" => Q := "010000";
         when x"4C2" => Q := "010000";
         when x"4C3" => Q := "010000";
         when x"4C4" => Q := "010000";
         when x"4C5" => Q := "010000";
         when x"4C6" => Q := "010000";
         when x"4C7" => Q := "011111";


-- CH=4D "M"
         when x"4D1" => Q := "010001";
         when x"4D2" => Q := "011011";
         when x"4D3" => Q := "010101";
         when x"4D4" => Q := "010101";
         when x"4D5" => Q := "010001";
         when x"4D6" => Q := "010001";
         when x"4D7" => Q := "010001";


-- CH=4E "N"
         when x"4E1" => Q := "010001";
         when x"4E2" => Q := "010001";
         when x"4E3" => Q := "011001";
         when x"4E4" => Q := "010101";
         when x"4E5" => Q := "010011";
         when x"4E6" => Q := "010001";
         when x"4E7" => Q := "010001";


-- CH=4F "O"
         when x"4F1" => Q := "001110";
         when x"4F2" => Q := "010001";
         when x"4F3" => Q := "010001";
         when x"4F4" => Q := "010001";
         when x"4F5" => Q := "010001";
         when x"4F6" => Q := "010001";
         when x"4F7" => Q := "001110";


-- CH=50 "P"
         when x"501" => Q := "011110";
         when x"502" => Q := "010001";
         when x"503" => Q := "010001";
         when x"504" => Q := "011110";
         when x"505" => Q := "010000";
         when x"506" => Q := "010000";
         when x"507" => Q := "010000";


-- CH=51 "Q"
         when x"511" => Q := "001110";
         when x"512" => Q := "010001";
         when x"513" => Q := "010001";
         when x"514" => Q := "010001";
         when x"515" => Q := "010101";
         when x"516" => Q := "010010";
         when x"517" => Q := "001101";


-- CH=52 "R"
         when x"521" => Q := "011110";
         when x"522" => Q := "010001";
         when x"523" => Q := "010001";
         when x"524" => Q := "011110";
         when x"525" => Q := "010100";
         when x"526" => Q := "010010";
         when x"527" => Q := "010001";


-- CH=53 "S"
         when x"531" => Q := "001110";
         when x"532" => Q := "010001";
         when x"533" => Q := "010000";
         when x"534" => Q := "001110";
         when x"535" => Q := "000001";
         when x"536" => Q := "010001";
         when x"537" => Q := "001110";


-- CH=54 "T"
         when x"541" => Q := "011111";
         when x"542" => Q := "000100";
         when x"543" => Q := "000100";
         when x"544" => Q := "000100";
         when x"545" => Q := "000100";
         when x"546" => Q := "000100";
         when x"547" => Q := "000100";


-- CH=55 "U"
         when x"551" => Q := "010001";
         when x"552" => Q := "010001";
         when x"553" => Q := "010001";
         when x"554" => Q := "010001";
         when x"555" => Q := "010001";
         when x"556" => Q := "010001";
         when x"557" => Q := "001110";


-- CH=56 "V"
         when x"561" => Q := "010001";
         when x"562" => Q := "010001";
         when x"563" => Q := "010001";
         when x"564" => Q := "001010";
         when x"565" => Q := "001010";
         when x"566" => Q := "000100";
         when x"567" => Q := "000100";


-- CH=57 "W"
         when x"571" => Q := "010001";
         when x"572" => Q := "010001";
         when x"573" => Q := "010001";
         when x"574" => Q := "010101";
         when x"575" => Q := "010101";
         when x"576" => Q := "010101";
         when x"577" => Q := "001010";


-- CH=58 "X"
         when x"581" => Q := "010001";
         when x"582" => Q := "010001";
         when x"583" => Q := "001010";
         when x"584" => Q := "000100";
         when x"585" => Q := "001010";
         when x"586" => Q := "010001";
         when x"587" => Q := "010001";


-- CH=59 "Y"
         when x"591" => Q := "010001";
         when x"592" => Q := "010001";
         when x"593" => Q := "001010";
         when x"594" => Q := "000100";
         when x"595" => Q := "000100";
         when x"596" => Q := "000100";
         when x"597" => Q := "000100";


-- CH=5A "Z"
         when x"5A1" => Q := "011111";
         when x"5A2" => Q := "000001";
         when x"5A3" => Q := "000010";
         when x"5A4" => Q := "000100";
         when x"5A5" => Q := "001000";
         when x"5A6" => Q := "010000";
         when x"5A7" => Q := "011111";


-- CH=5B "["
         when x"5B2" => Q := "000100";
         when x"5B3" => Q := "001000";
         when x"5B4" => Q := "011111";
         when x"5B5" => Q := "001000";
         when x"5B6" => Q := "000100";


-- CH=5C "\"
         when x"5C1" => Q := "010000";
         when x"5C2" => Q := "010000";
         when x"5C3" => Q := "010000";
         when x"5C4" => Q := "010000";
         when x"5C5" => Q := "010110";
         when x"5C6" => Q := "000001";
         when x"5C7" => Q := "000010";
         when x"5C8" => Q := "000100";
         when x"5C9" => Q := "000111";


-- CH=5D "]"
         when x"5D2" => Q := "000100";
         when x"5D3" => Q := "000010";
         when x"5D4" => Q := "011111";
         when x"5D5" => Q := "000010";
         when x"5D6" => Q := "000100";


-- CH=5E "^"
         when x"5E2" => Q := "000100";
         when x"5E3" => Q := "001110";
         when x"5E4" => Q := "010101";
         when x"5E5" => Q := "000100";
         when x"5E6" => Q := "000100";


-- CH=5F "_"
         when x"5F1" => Q := "001010";
         when x"5F2" => Q := "001010";
         when x"5F3" => Q := "011111";
         when x"5F4" => Q := "001010";
         when x"5F5" => Q := "011111";
         when x"5F6" => Q := "001010";
         when x"5F7" => Q := "001010";


-- CH=60 "`"
         when x"604" => Q := "011111";


-- CH=61 "a"
         when x"613" => Q := "001110";
         when x"614" => Q := "000001";
         when x"615" => Q := "001111";
         when x"616" => Q := "010001";
         when x"617" => Q := "001111";


-- CH=62 "b"
         when x"621" => Q := "010000";
         when x"622" => Q := "010000";
         when x"623" => Q := "011110";
         when x"624" => Q := "010001";
         when x"625" => Q := "010001";
         when x"626" => Q := "010001";
         when x"627" => Q := "011110";


-- CH=63 "c"
         when x"633" => Q := "001111";
         when x"634" => Q := "010000";
         when x"635" => Q := "010000";
         when x"636" => Q := "010000";
         when x"637" => Q := "001111";


-- CH=64 "d"
         when x"641" => Q := "000001";
         when x"642" => Q := "000001";
         when x"643" => Q := "001111";
         when x"644" => Q := "010001";
         when x"645" => Q := "010001";
         when x"646" => Q := "010001";
         when x"647" => Q := "001111";


-- CH=65 "e"
         when x"653" => Q := "001110";
         when x"654" => Q := "010001";
         when x"655" => Q := "011111";
         when x"656" => Q := "010000";
         when x"657" => Q := "001110";


-- CH=66 "f"
         when x"661" => Q := "000010";
         when x"662" => Q := "000100";
         when x"663" => Q := "000100";
         when x"664" => Q := "001110";
         when x"665" => Q := "000100";
         when x"666" => Q := "000100";
         when x"667" => Q := "000100";


-- CH=67 "g"
         when x"673" => Q := "001111";
         when x"674" => Q := "010001";
         when x"675" => Q := "010001";
         when x"676" => Q := "010001";
         when x"677" => Q := "001111";
         when x"678" => Q := "000001";
         when x"679" => Q := "001110";


-- CH=68 "h"
         when x"681" => Q := "010000";
         when x"682" => Q := "010000";
         when x"683" => Q := "011110";
         when x"684" => Q := "010001";
         when x"685" => Q := "010001";
         when x"686" => Q := "010001";
         when x"687" => Q := "010001";


-- CH=69 "i"
         when x"691" => Q := "000100";
         when x"693" => Q := "001100";
         when x"694" => Q := "000100";
         when x"695" => Q := "000100";
         when x"696" => Q := "000100";
         when x"697" => Q := "001110";


-- CH=6A "j"
         when x"6A1" => Q := "000100";
         when x"6A3" => Q := "000100";
         when x"6A4" => Q := "000100";
         when x"6A5" => Q := "000100";
         when x"6A6" => Q := "000100";
         when x"6A7" => Q := "000100";
         when x"6A8" => Q := "000100";
         when x"6A9" => Q := "001000";


-- CH=6B "k"
         when x"6B1" => Q := "001000";
         when x"6B2" => Q := "001000";
         when x"6B3" => Q := "001001";
         when x"6B4" => Q := "001010";
         when x"6B5" => Q := "001100";
         when x"6B6" => Q := "001010";
         when x"6B7" => Q := "001001";


-- CH=6C "l"
         when x"6C1" => Q := "001100";
         when x"6C2" => Q := "000100";
         when x"6C3" => Q := "000100";
         when x"6C4" => Q := "000100";
         when x"6C5" => Q := "000100";
         when x"6C6" => Q := "000100";
         when x"6C7" => Q := "001110";


-- CH=6D "m"
         when x"6D3" => Q := "011010";
         when x"6D4" => Q := "010101";
         when x"6D5" => Q := "010101";
         when x"6D6" => Q := "010101";
         when x"6D7" => Q := "010101";


-- CH=6E "n"
         when x"6E3" => Q := "011110";
         when x"6E4" => Q := "010001";
         when x"6E5" => Q := "010001";
         when x"6E6" => Q := "010001";
         when x"6E7" => Q := "010001";


-- CH=6F "o"
         when x"6F3" => Q := "001110";
         when x"6F4" => Q := "010001";
         when x"6F5" => Q := "010001";
         when x"6F6" => Q := "010001";
         when x"6F7" => Q := "001110";


-- CH=70 "p"
         when x"703" => Q := "011110";
         when x"704" => Q := "010001";
         when x"705" => Q := "010001";
         when x"706" => Q := "010001";
         when x"707" => Q := "011110";
         when x"708" => Q := "010000";
         when x"709" => Q := "010000";


-- CH=71 "q"
         when x"713" => Q := "001111";
         when x"714" => Q := "010001";
         when x"715" => Q := "010001";
         when x"716" => Q := "010001";
         when x"717" => Q := "001111";
         when x"718" => Q := "000001";
         when x"719" => Q := "000001";


-- CH=72 "r"
         when x"723" => Q := "001011";
         when x"724" => Q := "001100";
         when x"725" => Q := "001000";
         when x"726" => Q := "001000";
         when x"727" => Q := "001000";


-- CH=73 "s"
         when x"733" => Q := "001111";
         when x"734" => Q := "010000";
         when x"735" => Q := "001110";
         when x"736" => Q := "000001";
         when x"737" => Q := "011110";


-- CH=74 "t"
         when x"741" => Q := "000100";
         when x"742" => Q := "000100";
         when x"743" => Q := "001110";
         when x"744" => Q := "000100";
         when x"745" => Q := "000100";
         when x"746" => Q := "000100";
         when x"747" => Q := "000010";


-- CH=75 "u"
         when x"753" => Q := "010001";
         when x"754" => Q := "010001";
         when x"755" => Q := "010001";
         when x"756" => Q := "010001";
         when x"757" => Q := "001111";


-- CH=76 "v"
         when x"763" => Q := "010001";
         when x"764" => Q := "010001";
         when x"765" => Q := "001010";
         when x"766" => Q := "001010";
         when x"767" => Q := "000100";


-- CH=77 "w"
         when x"773" => Q := "010001";
         when x"774" => Q := "010001";
         when x"775" => Q := "010101";
         when x"776" => Q := "010101";
         when x"777" => Q := "001010";


-- CH=78 "x"
         when x"783" => Q := "010001";
         when x"784" => Q := "001010";
         when x"785" => Q := "000100";
         when x"786" => Q := "001010";
         when x"787" => Q := "010001";


-- CH=79 "y"
         when x"793" => Q := "010001";
         when x"794" => Q := "010001";
         when x"795" => Q := "010001";
         when x"796" => Q := "010001";
         when x"797" => Q := "001111";
         when x"798" => Q := "000001";
         when x"799" => Q := "001110";


-- CH=7A "z"
         when x"7A3" => Q := "011111";
         when x"7A4" => Q := "000010";
         when x"7A5" => Q := "000100";
         when x"7A6" => Q := "001000";
         when x"7A7" => Q := "011111";


-- CH=7B "{"
         when x"7B1" => Q := "001000";
         when x"7B2" => Q := "001000";
         when x"7B3" => Q := "001000";
         when x"7B4" => Q := "001000";
         when x"7B5" => Q := "001001";
         when x"7B6" => Q := "000011";
         when x"7B7" => Q := "000101";
         when x"7B8" => Q := "000111";
         when x"7B9" => Q := "000001";


-- CH=7C "|"
         when x"7C1" => Q := "001010";
         when x"7C2" => Q := "001010";
         when x"7C3" => Q := "001010";
         when x"7C4" => Q := "001010";
         when x"7C5" => Q := "001010";
         when x"7C6" => Q := "001010";
         when x"7C7" => Q := "001010";


-- CH=7D "}"
         when x"7D1" => Q := "011000";
         when x"7D2" => Q := "000100";
         when x"7D3" => Q := "011000";
         when x"7D4" => Q := "000100";
         when x"7D5" => Q := "011001";
         when x"7D6" => Q := "000011";
         when x"7D7" => Q := "000101";
         when x"7D8" => Q := "000111";
         when x"7D9" => Q := "000001";


-- CH=7E "~"
         when x"7E2" => Q := "000100";
         when x"7E4" => Q := "011111";
         when x"7E6" => Q := "000100";


-- CH=7F ""
         when x"7F1" => Q := "011111";
         when x"7F2" => Q := "011111";
         when x"7F3" => Q := "011111";
         when x"7F4" => Q := "011111";
         when x"7F5" => Q := "011111";
         when x"7F6" => Q := "011111";
         when x"7F7" => Q := "011111";

	   	when others => Q := (others => '0');

	   end case;

	   if A(11) = '1' and A(9) = '1' then
         case to_integer(unsigned(A(3 downto 0))) is
            when 0|1|2 =>
               Q := A(4) & A(4) & A(4) & A(5) & A(5) & A(5);
            when 3|4|5|6 =>
               Q := A(6) & A(6) & A(6) & A(7) & A(7) & A(7);
            when others =>
               Q := A(8) & A(8) & A(8) & A(10) & A(10) & A(10);
         end case;
         if r_switch = '0' then
            QA <= "10" & Q;
         else
            QB <= "10" & Q;
         end if;
      else
           -- text / blast
    	   if r_switch = '0' then
    	   	QA <= "00" & Q;
    	   else
    	   	QB <= "00" & Q;
    	   end if;
      end if;

		r_switch <= not r_switch;
	end if;

end process;

end RTL;