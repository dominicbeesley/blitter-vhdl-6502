-- hdmi_serial.vhd

-- Generated using ACDS version 20.1 720

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity hdmi_serial is
	port (
		tx_inclock   : in  std_logic                     := '0';             --   tx_inclock.tx_inclock
		tx_syncclock : in  std_logic                     := '0';             -- tx_syncclock.tx_syncclock
		tx_in        : in  std_logic_vector(39 downto 0) := (others => '0'); --        tx_in.tx_in
		tx_out       : out std_logic_vector(3 downto 0)                      --       tx_out.tx_out
	);
end entity hdmi_serial;

architecture rtl of hdmi_serial is
	component altera_soft_lvds_tx_SzWJL is
		port (
			tx_inclock   : in  std_logic                     := 'X';             -- tx_inclock
			tx_syncclock : in  std_logic                     := 'X';             -- tx_syncclock
			tx_in        : in  std_logic_vector(39 downto 0) := (others => 'X'); -- tx_in
			tx_out       : out std_logic_vector(3 downto 0);                     -- tx_out
			tx_outclock  : out std_logic;                                        -- tx_outclock
			tx_coreclock : out std_logic;                                        -- tx_coreclock
			tx_locked    : out std_logic                                         -- tx_locked
		);
	end component altera_soft_lvds_tx_SzWJL;

begin

	hdmi_serial_inst : component altera_soft_lvds_tx_SzWJL
		port map (
			tx_inclock   => tx_inclock,   --   tx_inclock.tx_inclock
			tx_syncclock => tx_syncclock, -- tx_syncclock.tx_syncclock
			tx_in        => tx_in,        --        tx_in.tx_in
			tx_out       => tx_out,       --       tx_out.tx_out
			tx_outclock  => open,         --  (terminated)
			tx_coreclock => open,         --  (terminated)
			tx_locked    => open          --  (terminated)
		);

end architecture rtl; -- of hdmi_serial
