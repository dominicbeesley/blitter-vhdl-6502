-- MIT License
-- -----------------------------------------------------------------------------
-- Copyright (c) 2021 Dominic Beesley https://github.com/dominicbeesley
--
-- Permission is hereby granted, free of charge, to any person obtaining a copy
-- of this software and associated documentation files (the "Software"), to deal
-- in the Software without restriction, including without limitation the rights
-- to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
-- copies of the Software, and to permit persons to whom the Software is
-- furnished to do so, subject to the following conditions:
--
-- The above copyright notice and this permission notice shall be included in
-- all copies or substantial portions of the Software.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
-- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
-- FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
-- AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
-- LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
-- OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
-- THE SOFTWARE.
-- ----------------------------------------------------------------------


-- Company: 				Dossytronics
-- Engineer: 				Dominic Beesley
-- 
-- Create Date:    		29/1/2022
-- Design Name: 
-- Module Name:    		work.real80188
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 			mimic the external behaviour of a 80188 CPU
-- Dependencies: 
--
-- Revision: 
-- Additional Comments: CAUTION: this is very much a work in progress and
--								only mimics the most basic parts of an 80188
--								
--
----------------------------------------------------------------------------------



library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity real80188_tb is
	generic (
		Tcico		:	time := 17 ns
	);
	port(

		X1_i		: in 	std_logic;

		CLKOUT_o	: out std_logic

	);
end real80188_tb;

architecture behavioral of real80188_tb is
	signal	r_CLK_int	: std_logic;
	signal	i_CLKOUT		: std_logic;
begin


	p_X1:process(X1_i)
	begin
		if falling_edge(X1_i) then
			if r_CLK_int = '0' then
				r_CLK_int <= '1';
			else
				r_CLK_int <= '0';
			end if;
		end if;
	end process;

	i_CLKOUT <= r_CLK_int after Tcico;
	CLKOUT_o <= i_CLKOUT;


end behavioral;