library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity saa5050_rom_dual_port is
    generic (
        ADDR_WIDTH       : integer := 12;
        DATA_WIDTH       : integer := 8
    );
    port(
        clock    : in  std_logic;
        addressA : in  std_logic_vector(11 downto 0);
        QA       : out std_logic_vector(7 downto 0);
        addressB : in  std_logic_vector(11 downto 0);
        QB       : out std_logic_vector(7 downto 0)
  );
end saa5050_rom_dual_port;

architecture RTL of saa5050_rom_dual_port is

signal	r_switch : std_logic := '0';

begin

p:process(CLOCK)
variable A:std_logic_vector(11 downto 0);
variable Q:std_logic_vector(5 downto 0);
variable TOP:std_logic;
begin

	if (rising_edge(CLOCK)) then
		if (r_switch = '0') then
			A := addressA;
		else
			A := addressB;
		end if;

		case (A) is

-- CH=21 "!"
         when x"211" => Q := "000100";
         when x"212" => Q := "000100";
         when x"213" => Q := "000100";
         when x"214" => Q := "000100";
         when x"215" => Q := "000100";
         when x"217" => Q := "000100";


-- CH=22 """
         when x"221" => Q := "001010";
         when x"222" => Q := "001010";
         when x"223" => Q := "001010";


-- CH=23 "#"
         when x"231" => Q := "000110";
         when x"232" => Q := "001001";
         when x"233" => Q := "001000";
         when x"234" => Q := "011100";
         when x"235" => Q := "001000";
         when x"236" => Q := "001000";
         when x"237" => Q := "011111";


-- CH=24 "$"
         when x"241" => Q := "001110";
         when x"242" => Q := "010101";
         when x"243" => Q := "010100";
         when x"244" => Q := "001110";
         when x"245" => Q := "000101";
         when x"246" => Q := "010101";
         when x"247" => Q := "001110";


-- CH=25 "%"
         when x"251" => Q := "011000";
         when x"252" => Q := "011001";
         when x"253" => Q := "000010";
         when x"254" => Q := "000100";
         when x"255" => Q := "001000";
         when x"256" => Q := "010011";
         when x"257" => Q := "000011";


-- CH=26 "&"
         when x"261" => Q := "001000";
         when x"262" => Q := "010100";
         when x"263" => Q := "010100";
         when x"264" => Q := "001000";
         when x"265" => Q := "010101";
         when x"266" => Q := "010010";
         when x"267" => Q := "001101";


-- CH=27 "'"
         when x"271" => Q := "000100";
         when x"272" => Q := "000100";
         when x"273" => Q := "000100";


-- CH=28 "("
         when x"281" => Q := "000010";
         when x"282" => Q := "000100";
         when x"283" => Q := "001000";
         when x"284" => Q := "001000";
         when x"285" => Q := "001000";
         when x"286" => Q := "000100";
         when x"287" => Q := "000010";


-- CH=29 ")"
         when x"291" => Q := "001000";
         when x"292" => Q := "000100";
         when x"293" => Q := "000010";
         when x"294" => Q := "000010";
         when x"295" => Q := "000010";
         when x"296" => Q := "000100";
         when x"297" => Q := "001000";


-- CH=2A "*"
         when x"2A1" => Q := "000100";
         when x"2A2" => Q := "010101";
         when x"2A3" => Q := "001110";
         when x"2A4" => Q := "000100";
         when x"2A5" => Q := "001110";
         when x"2A6" => Q := "010101";
         when x"2A7" => Q := "000100";


-- CH=2B "+"
         when x"2B2" => Q := "000100";
         when x"2B3" => Q := "000100";
         when x"2B4" => Q := "011111";
         when x"2B5" => Q := "000100";
         when x"2B6" => Q := "000100";


-- CH=2C ","
         when x"2C6" => Q := "000100";
         when x"2C7" => Q := "000100";
         when x"2C8" => Q := "001000";


-- CH=2D "-"
         when x"2D4" => Q := "001110";


-- CH=2E "."
         when x"2E7" => Q := "000100";


-- CH=2F "/"
         when x"2F2" => Q := "000001";
         when x"2F3" => Q := "000010";
         when x"2F4" => Q := "000100";
         when x"2F5" => Q := "001000";
         when x"2F6" => Q := "010000";


-- CH=30 "0"
         when x"301" => Q := "000100";
         when x"302" => Q := "001010";
         when x"303" => Q := "010001";
         when x"304" => Q := "010001";
         when x"305" => Q := "010001";
         when x"306" => Q := "001010";
         when x"307" => Q := "000100";


-- CH=31 "1"
         when x"311" => Q := "000100";
         when x"312" => Q := "001100";
         when x"313" => Q := "000100";
         when x"314" => Q := "000100";
         when x"315" => Q := "000100";
         when x"316" => Q := "000100";
         when x"317" => Q := "001110";


-- CH=32 "2"
         when x"321" => Q := "001110";
         when x"322" => Q := "010001";
         when x"323" => Q := "000001";
         when x"324" => Q := "000110";
         when x"325" => Q := "001000";
         when x"326" => Q := "010000";
         when x"327" => Q := "011111";


-- CH=33 "3"
         when x"331" => Q := "011111";
         when x"332" => Q := "000001";
         when x"333" => Q := "000010";
         when x"334" => Q := "000110";
         when x"335" => Q := "000001";
         when x"336" => Q := "010001";
         when x"337" => Q := "001110";


-- CH=34 "4"
         when x"341" => Q := "000010";
         when x"342" => Q := "000110";
         when x"343" => Q := "001010";
         when x"344" => Q := "010010";
         when x"345" => Q := "011111";
         when x"346" => Q := "000010";
         when x"347" => Q := "000010";


-- CH=35 "5"
         when x"351" => Q := "011111";
         when x"352" => Q := "010000";
         when x"353" => Q := "011110";
         when x"354" => Q := "000001";
         when x"355" => Q := "000001";
         when x"356" => Q := "010001";
         when x"357" => Q := "001110";


-- CH=36 "6"
         when x"361" => Q := "000110";
         when x"362" => Q := "001000";
         when x"363" => Q := "010000";
         when x"364" => Q := "011110";
         when x"365" => Q := "010001";
         when x"366" => Q := "010001";
         when x"367" => Q := "001110";


-- CH=37 "7"
         when x"371" => Q := "011111";
         when x"372" => Q := "000001";
         when x"373" => Q := "000010";
         when x"374" => Q := "000100";
         when x"375" => Q := "001000";
         when x"376" => Q := "001000";
         when x"377" => Q := "001000";


-- CH=38 "8"
         when x"381" => Q := "001110";
         when x"382" => Q := "010001";
         when x"383" => Q := "010001";
         when x"384" => Q := "001110";
         when x"385" => Q := "010001";
         when x"386" => Q := "010001";
         when x"387" => Q := "001110";


-- CH=39 "9"
         when x"391" => Q := "001110";
         when x"392" => Q := "010001";
         when x"393" => Q := "010001";
         when x"394" => Q := "001111";
         when x"395" => Q := "000001";
         when x"396" => Q := "000010";
         when x"397" => Q := "001100";


-- CH=3A ":"
         when x"3A3" => Q := "000100";
         when x"3A7" => Q := "000100";


-- CH=3B ";"
         when x"3B3" => Q := "000100";
         when x"3B6" => Q := "000100";
         when x"3B7" => Q := "000100";
         when x"3B8" => Q := "001000";


-- CH=3C "<"
         when x"3C1" => Q := "000010";
         when x"3C2" => Q := "000100";
         when x"3C3" => Q := "001000";
         when x"3C4" => Q := "010000";
         when x"3C5" => Q := "001000";
         when x"3C6" => Q := "000100";
         when x"3C7" => Q := "000010";


-- CH=3D "="
         when x"3D3" => Q := "011111";
         when x"3D5" => Q := "011111";


-- CH=3E ">"
         when x"3E1" => Q := "001000";
         when x"3E2" => Q := "000100";
         when x"3E3" => Q := "000010";
         when x"3E4" => Q := "000001";
         when x"3E5" => Q := "000010";
         when x"3E6" => Q := "000100";
         when x"3E7" => Q := "001000";


-- CH=3F "?"
         when x"3F1" => Q := "001110";
         when x"3F2" => Q := "010001";
         when x"3F3" => Q := "000010";
         when x"3F4" => Q := "000100";
         when x"3F5" => Q := "000100";
         when x"3F7" => Q := "000100";


-- CH=40 "@"
         when x"401" => Q := "001110";
         when x"402" => Q := "010001";
         when x"403" => Q := "010111";
         when x"404" => Q := "010101";
         when x"405" => Q := "010111";
         when x"406" => Q := "010000";
         when x"407" => Q := "001110";


-- CH=41 "A"
         when x"411" => Q := "000100";
         when x"412" => Q := "001010";
         when x"413" => Q := "010001";
         when x"414" => Q := "010001";
         when x"415" => Q := "011111";
         when x"416" => Q := "010001";
         when x"417" => Q := "010001";


-- CH=42 "B"
         when x"421" => Q := "011110";
         when x"422" => Q := "010001";
         when x"423" => Q := "010001";
         when x"424" => Q := "011110";
         when x"425" => Q := "010001";
         when x"426" => Q := "010001";
         when x"427" => Q := "011110";


-- CH=43 "C"
         when x"431" => Q := "001110";
         when x"432" => Q := "010001";
         when x"433" => Q := "010000";
         when x"434" => Q := "010000";
         when x"435" => Q := "010000";
         when x"436" => Q := "010001";
         when x"437" => Q := "001110";


-- CH=44 "D"
         when x"441" => Q := "011110";
         when x"442" => Q := "010001";
         when x"443" => Q := "010001";
         when x"444" => Q := "010001";
         when x"445" => Q := "010001";
         when x"446" => Q := "010001";
         when x"447" => Q := "011110";


-- CH=45 "E"
         when x"451" => Q := "011111";
         when x"452" => Q := "010000";
         when x"453" => Q := "010000";
         when x"454" => Q := "011110";
         when x"455" => Q := "010000";
         when x"456" => Q := "010000";
         when x"457" => Q := "011111";


-- CH=46 "F"
         when x"461" => Q := "011111";
         when x"462" => Q := "010000";
         when x"463" => Q := "010000";
         when x"464" => Q := "011110";
         when x"465" => Q := "010000";
         when x"466" => Q := "010000";
         when x"467" => Q := "010000";


-- CH=47 "G"
         when x"471" => Q := "001110";
         when x"472" => Q := "010001";
         when x"473" => Q := "010000";
         when x"474" => Q := "010000";
         when x"475" => Q := "010011";
         when x"476" => Q := "010001";
         when x"477" => Q := "001111";


-- CH=48 "H"
         when x"481" => Q := "010001";
         when x"482" => Q := "010001";
         when x"483" => Q := "010001";
         when x"484" => Q := "011111";
         when x"485" => Q := "010001";
         when x"486" => Q := "010001";
         when x"487" => Q := "010001";


-- CH=49 "I"
         when x"491" => Q := "001110";
         when x"492" => Q := "000100";
         when x"493" => Q := "000100";
         when x"494" => Q := "000100";
         when x"495" => Q := "000100";
         when x"496" => Q := "000100";
         when x"497" => Q := "001110";


-- CH=4A "J"
         when x"4A1" => Q := "000001";
         when x"4A2" => Q := "000001";
         when x"4A3" => Q := "000001";
         when x"4A4" => Q := "000001";
         when x"4A5" => Q := "000001";
         when x"4A6" => Q := "010001";
         when x"4A7" => Q := "001110";


-- CH=4B "K"
         when x"4B1" => Q := "010001";
         when x"4B2" => Q := "010010";
         when x"4B3" => Q := "010100";
         when x"4B4" => Q := "011000";
         when x"4B5" => Q := "010100";
         when x"4B6" => Q := "010010";
         when x"4B7" => Q := "010001";


-- CH=4C "L"
         when x"4C1" => Q := "010000";
         when x"4C2" => Q := "010000";
         when x"4C3" => Q := "010000";
         when x"4C4" => Q := "010000";
         when x"4C5" => Q := "010000";
         when x"4C6" => Q := "010000";
         when x"4C7" => Q := "011111";


-- CH=4D "M"
         when x"4D1" => Q := "010001";
         when x"4D2" => Q := "011011";
         when x"4D3" => Q := "010101";
         when x"4D4" => Q := "010101";
         when x"4D5" => Q := "010001";
         when x"4D6" => Q := "010001";
         when x"4D7" => Q := "010001";


-- CH=4E "N"
         when x"4E1" => Q := "010001";
         when x"4E2" => Q := "010001";
         when x"4E3" => Q := "011001";
         when x"4E4" => Q := "010101";
         when x"4E5" => Q := "010011";
         when x"4E6" => Q := "010001";
         when x"4E7" => Q := "010001";


-- CH=4F "O"
         when x"4F1" => Q := "001110";
         when x"4F2" => Q := "010001";
         when x"4F3" => Q := "010001";
         when x"4F4" => Q := "010001";
         when x"4F5" => Q := "010001";
         when x"4F6" => Q := "010001";
         when x"4F7" => Q := "001110";


-- CH=50 "P"
         when x"501" => Q := "011110";
         when x"502" => Q := "010001";
         when x"503" => Q := "010001";
         when x"504" => Q := "011110";
         when x"505" => Q := "010000";
         when x"506" => Q := "010000";
         when x"507" => Q := "010000";


-- CH=51 "Q"
         when x"511" => Q := "001110";
         when x"512" => Q := "010001";
         when x"513" => Q := "010001";
         when x"514" => Q := "010001";
         when x"515" => Q := "010101";
         when x"516" => Q := "010010";
         when x"517" => Q := "001101";


-- CH=52 "R"
         when x"521" => Q := "011110";
         when x"522" => Q := "010001";
         when x"523" => Q := "010001";
         when x"524" => Q := "011110";
         when x"525" => Q := "010100";
         when x"526" => Q := "010010";
         when x"527" => Q := "010001";


-- CH=53 "S"
         when x"531" => Q := "001110";
         when x"532" => Q := "010001";
         when x"533" => Q := "010000";
         when x"534" => Q := "001110";
         when x"535" => Q := "000001";
         when x"536" => Q := "010001";
         when x"537" => Q := "001110";


-- CH=54 "T"
         when x"541" => Q := "011111";
         when x"542" => Q := "000100";
         when x"543" => Q := "000100";
         when x"544" => Q := "000100";
         when x"545" => Q := "000100";
         when x"546" => Q := "000100";
         when x"547" => Q := "000100";


-- CH=55 "U"
         when x"551" => Q := "010001";
         when x"552" => Q := "010001";
         when x"553" => Q := "010001";
         when x"554" => Q := "010001";
         when x"555" => Q := "010001";
         when x"556" => Q := "010001";
         when x"557" => Q := "001110";


-- CH=56 "V"
         when x"561" => Q := "010001";
         when x"562" => Q := "010001";
         when x"563" => Q := "010001";
         when x"564" => Q := "001010";
         when x"565" => Q := "001010";
         when x"566" => Q := "000100";
         when x"567" => Q := "000100";


-- CH=57 "W"
         when x"571" => Q := "010001";
         when x"572" => Q := "010001";
         when x"573" => Q := "010001";
         when x"574" => Q := "010101";
         when x"575" => Q := "010101";
         when x"576" => Q := "010101";
         when x"577" => Q := "001010";


-- CH=58 "X"
         when x"581" => Q := "010001";
         when x"582" => Q := "010001";
         when x"583" => Q := "001010";
         when x"584" => Q := "000100";
         when x"585" => Q := "001010";
         when x"586" => Q := "010001";
         when x"587" => Q := "010001";


-- CH=59 "Y"
         when x"591" => Q := "010001";
         when x"592" => Q := "010001";
         when x"593" => Q := "001010";
         when x"594" => Q := "000100";
         when x"595" => Q := "000100";
         when x"596" => Q := "000100";
         when x"597" => Q := "000100";


-- CH=5A "Z"
         when x"5A1" => Q := "011111";
         when x"5A2" => Q := "000001";
         when x"5A3" => Q := "000010";
         when x"5A4" => Q := "000100";
         when x"5A5" => Q := "001000";
         when x"5A6" => Q := "010000";
         when x"5A7" => Q := "011111";


-- CH=5B "["
         when x"5B2" => Q := "000100";
         when x"5B3" => Q := "001000";
         when x"5B4" => Q := "011111";
         when x"5B5" => Q := "001000";
         when x"5B6" => Q := "000100";


-- CH=5C "\"
         when x"5C1" => Q := "010000";
         when x"5C2" => Q := "010000";
         when x"5C3" => Q := "010000";
         when x"5C4" => Q := "010000";
         when x"5C5" => Q := "010110";
         when x"5C6" => Q := "000001";
         when x"5C7" => Q := "000010";
         when x"5C8" => Q := "000100";
         when x"5C9" => Q := "000111";


-- CH=5D "]"
         when x"5D2" => Q := "000100";
         when x"5D3" => Q := "000010";
         when x"5D4" => Q := "011111";
         when x"5D5" => Q := "000010";
         when x"5D6" => Q := "000100";


-- CH=5E "^"
         when x"5E2" => Q := "000100";
         when x"5E3" => Q := "001110";
         when x"5E4" => Q := "010101";
         when x"5E5" => Q := "000100";
         when x"5E6" => Q := "000100";


-- CH=5F "_"
         when x"5F1" => Q := "001010";
         when x"5F2" => Q := "001010";
         when x"5F3" => Q := "011111";
         when x"5F4" => Q := "001010";
         when x"5F5" => Q := "011111";
         when x"5F6" => Q := "001010";
         when x"5F7" => Q := "001010";


-- CH=60 "`"
         when x"604" => Q := "011111";


-- CH=61 "a"
         when x"613" => Q := "001110";
         when x"614" => Q := "000001";
         when x"615" => Q := "001111";
         when x"616" => Q := "010001";
         when x"617" => Q := "001111";


-- CH=62 "b"
         when x"621" => Q := "010000";
         when x"622" => Q := "010000";
         when x"623" => Q := "011110";
         when x"624" => Q := "010001";
         when x"625" => Q := "010001";
         when x"626" => Q := "010001";
         when x"627" => Q := "011110";


-- CH=63 "c"
         when x"633" => Q := "001111";
         when x"634" => Q := "010000";
         when x"635" => Q := "010000";
         when x"636" => Q := "010000";
         when x"637" => Q := "001111";


-- CH=64 "d"
         when x"641" => Q := "000001";
         when x"642" => Q := "000001";
         when x"643" => Q := "001111";
         when x"644" => Q := "010001";
         when x"645" => Q := "010001";
         when x"646" => Q := "010001";
         when x"647" => Q := "001111";


-- CH=65 "e"
         when x"653" => Q := "001110";
         when x"654" => Q := "010001";
         when x"655" => Q := "011111";
         when x"656" => Q := "010000";
         when x"657" => Q := "001110";


-- CH=66 "f"
         when x"661" => Q := "000010";
         when x"662" => Q := "000100";
         when x"663" => Q := "000100";
         when x"664" => Q := "001110";
         when x"665" => Q := "000100";
         when x"666" => Q := "000100";
         when x"667" => Q := "000100";


-- CH=67 "g"
         when x"673" => Q := "001111";
         when x"674" => Q := "010001";
         when x"675" => Q := "010001";
         when x"676" => Q := "010001";
         when x"677" => Q := "001111";
         when x"678" => Q := "000001";
         when x"679" => Q := "001110";


-- CH=68 "h"
         when x"681" => Q := "010000";
         when x"682" => Q := "010000";
         when x"683" => Q := "011110";
         when x"684" => Q := "010001";
         when x"685" => Q := "010001";
         when x"686" => Q := "010001";
         when x"687" => Q := "010001";


-- CH=69 "i"
         when x"691" => Q := "000100";
         when x"693" => Q := "001100";
         when x"694" => Q := "000100";
         when x"695" => Q := "000100";
         when x"696" => Q := "000100";
         when x"697" => Q := "001110";


-- CH=6A "j"
         when x"6A1" => Q := "000100";
         when x"6A3" => Q := "000100";
         when x"6A4" => Q := "000100";
         when x"6A5" => Q := "000100";
         when x"6A6" => Q := "000100";
         when x"6A7" => Q := "000100";
         when x"6A8" => Q := "000100";
         when x"6A9" => Q := "001000";


-- CH=6B "k"
         when x"6B1" => Q := "001000";
         when x"6B2" => Q := "001000";
         when x"6B3" => Q := "001001";
         when x"6B4" => Q := "001010";
         when x"6B5" => Q := "001100";
         when x"6B6" => Q := "001010";
         when x"6B7" => Q := "001001";


-- CH=6C "l"
         when x"6C1" => Q := "001100";
         when x"6C2" => Q := "000100";
         when x"6C3" => Q := "000100";
         when x"6C4" => Q := "000100";
         when x"6C5" => Q := "000100";
         when x"6C6" => Q := "000100";
         when x"6C7" => Q := "001110";


-- CH=6D "m"
         when x"6D3" => Q := "011010";
         when x"6D4" => Q := "010101";
         when x"6D5" => Q := "010101";
         when x"6D6" => Q := "010101";
         when x"6D7" => Q := "010101";


-- CH=6E "n"
         when x"6E3" => Q := "011110";
         when x"6E4" => Q := "010001";
         when x"6E5" => Q := "010001";
         when x"6E6" => Q := "010001";
         when x"6E7" => Q := "010001";


-- CH=6F "o"
         when x"6F3" => Q := "001110";
         when x"6F4" => Q := "010001";
         when x"6F5" => Q := "010001";
         when x"6F6" => Q := "010001";
         when x"6F7" => Q := "001110";


-- CH=70 "p"
         when x"703" => Q := "011110";
         when x"704" => Q := "010001";
         when x"705" => Q := "010001";
         when x"706" => Q := "010001";
         when x"707" => Q := "011110";
         when x"708" => Q := "010000";
         when x"709" => Q := "010000";


-- CH=71 "q"
         when x"713" => Q := "001111";
         when x"714" => Q := "010001";
         when x"715" => Q := "010001";
         when x"716" => Q := "010001";
         when x"717" => Q := "001111";
         when x"718" => Q := "000001";
         when x"719" => Q := "000001";


-- CH=72 "r"
         when x"723" => Q := "001011";
         when x"724" => Q := "001100";
         when x"725" => Q := "001000";
         when x"726" => Q := "001000";
         when x"727" => Q := "001000";


-- CH=73 "s"
         when x"733" => Q := "001111";
         when x"734" => Q := "010000";
         when x"735" => Q := "001110";
         when x"736" => Q := "000001";
         when x"737" => Q := "011110";


-- CH=74 "t"
         when x"741" => Q := "000100";
         when x"742" => Q := "000100";
         when x"743" => Q := "001110";
         when x"744" => Q := "000100";
         when x"745" => Q := "000100";
         when x"746" => Q := "000100";
         when x"747" => Q := "000010";


-- CH=75 "u"
         when x"753" => Q := "010001";
         when x"754" => Q := "010001";
         when x"755" => Q := "010001";
         when x"756" => Q := "010001";
         when x"757" => Q := "001111";


-- CH=76 "v"
         when x"763" => Q := "010001";
         when x"764" => Q := "010001";
         when x"765" => Q := "001010";
         when x"766" => Q := "001010";
         when x"767" => Q := "000100";


-- CH=77 "w"
         when x"773" => Q := "010001";
         when x"774" => Q := "010001";
         when x"775" => Q := "010101";
         when x"776" => Q := "010101";
         when x"777" => Q := "001010";


-- CH=78 "x"
         when x"783" => Q := "010001";
         when x"784" => Q := "001010";
         when x"785" => Q := "000100";
         when x"786" => Q := "001010";
         when x"787" => Q := "010001";


-- CH=79 "y"
         when x"793" => Q := "010001";
         when x"794" => Q := "010001";
         when x"795" => Q := "010001";
         when x"796" => Q := "010001";
         when x"797" => Q := "001111";
         when x"798" => Q := "000001";
         when x"799" => Q := "001110";


-- CH=7A "z"
         when x"7A3" => Q := "011111";
         when x"7A4" => Q := "000010";
         when x"7A5" => Q := "000100";
         when x"7A6" => Q := "001000";
         when x"7A7" => Q := "011111";


-- CH=7B "{"
         when x"7B1" => Q := "001000";
         when x"7B2" => Q := "001000";
         when x"7B3" => Q := "001000";
         when x"7B4" => Q := "001000";
         when x"7B5" => Q := "001001";
         when x"7B6" => Q := "000011";
         when x"7B7" => Q := "000101";
         when x"7B8" => Q := "000111";
         when x"7B9" => Q := "000001";


-- CH=7C "|"
         when x"7C1" => Q := "001010";
         when x"7C2" => Q := "001010";
         when x"7C3" => Q := "001010";
         when x"7C4" => Q := "001010";
         when x"7C5" => Q := "001010";
         when x"7C6" => Q := "001010";
         when x"7C7" => Q := "001010";


-- CH=7D "}"
         when x"7D1" => Q := "011000";
         when x"7D2" => Q := "000100";
         when x"7D3" => Q := "011000";
         when x"7D4" => Q := "000100";
         when x"7D5" => Q := "011001";
         when x"7D6" => Q := "000011";
         when x"7D7" => Q := "000101";
         when x"7D8" => Q := "000111";
         when x"7D9" => Q := "000001";


-- CH=7E "~"
         when x"7E2" => Q := "000100";
         when x"7E4" => Q := "011111";
         when x"7E6" => Q := "000100";


-- CH=7F ""
         when x"7F1" => Q := "011111";
         when x"7F2" => Q := "011111";
         when x"7F3" => Q := "011111";
         when x"7F4" => Q := "011111";
         when x"7F5" => Q := "011111";
         when x"7F6" => Q := "011111";
         when x"7F7" => Q := "011111";


-- CH=A1 
         when x"A10" => Q := "111000";
         when x"A11" => Q := "111000";
         when x"A12" => Q := "111000";


-- CH=A2 
         when x"A20" => Q := "000111";
         when x"A21" => Q := "000111";
         when x"A22" => Q := "000111";


-- CH=A3 
         when x"A30" => Q := "111111";
         when x"A31" => Q := "111111";
         when x"A32" => Q := "111111";


-- CH=A4 
         when x"A43" => Q := "111000";
         when x"A44" => Q := "111000";
         when x"A45" => Q := "111000";
         when x"A46" => Q := "111000";


-- CH=A5 
         when x"A50" => Q := "111000";
         when x"A51" => Q := "111000";
         when x"A52" => Q := "111000";
         when x"A53" => Q := "111000";
         when x"A54" => Q := "111000";
         when x"A55" => Q := "111000";
         when x"A56" => Q := "111000";


-- CH=A6 
         when x"A60" => Q := "000111";
         when x"A61" => Q := "000111";
         when x"A62" => Q := "000111";
         when x"A63" => Q := "111000";
         when x"A64" => Q := "111000";
         when x"A65" => Q := "111000";
         when x"A66" => Q := "111000";


-- CH=A7 
         when x"A70" => Q := "111111";
         when x"A71" => Q := "111111";
         when x"A72" => Q := "111111";
         when x"A73" => Q := "111000";
         when x"A74" => Q := "111000";
         when x"A75" => Q := "111000";
         when x"A76" => Q := "111000";


-- CH=A8 
         when x"A83" => Q := "000111";
         when x"A84" => Q := "000111";
         when x"A85" => Q := "000111";
         when x"A86" => Q := "000111";


-- CH=A9 
         when x"A90" => Q := "111000";
         when x"A91" => Q := "111000";
         when x"A92" => Q := "111000";
         when x"A93" => Q := "000111";
         when x"A94" => Q := "000111";
         when x"A95" => Q := "000111";
         when x"A96" => Q := "000111";


-- CH=AA 
         when x"AA0" => Q := "000111";
         when x"AA1" => Q := "000111";
         when x"AA2" => Q := "000111";
         when x"AA3" => Q := "000111";
         when x"AA4" => Q := "000111";
         when x"AA5" => Q := "000111";
         when x"AA6" => Q := "000111";


-- CH=AB 
         when x"AB0" => Q := "111111";
         when x"AB1" => Q := "111111";
         when x"AB2" => Q := "111111";
         when x"AB3" => Q := "000111";
         when x"AB4" => Q := "000111";
         when x"AB5" => Q := "000111";
         when x"AB6" => Q := "000111";


-- CH=AC 
         when x"AC3" => Q := "111111";
         when x"AC4" => Q := "111111";
         when x"AC5" => Q := "111111";
         when x"AC6" => Q := "111111";


-- CH=AD 
         when x"AD0" => Q := "111000";
         when x"AD1" => Q := "111000";
         when x"AD2" => Q := "111000";
         when x"AD3" => Q := "111111";
         when x"AD4" => Q := "111111";
         when x"AD5" => Q := "111111";
         when x"AD6" => Q := "111111";


-- CH=AE 
         when x"AE0" => Q := "000111";
         when x"AE1" => Q := "000111";
         when x"AE2" => Q := "000111";
         when x"AE3" => Q := "111111";
         when x"AE4" => Q := "111111";
         when x"AE5" => Q := "111111";
         when x"AE6" => Q := "111111";


-- CH=AF 
         when x"AF0" => Q := "111111";
         when x"AF1" => Q := "111111";
         when x"AF2" => Q := "111111";
         when x"AF3" => Q := "111111";
         when x"AF4" => Q := "111111";
         when x"AF5" => Q := "111111";
         when x"AF6" => Q := "111111";


-- CH=B0 
         when x"B07" => Q := "111000";
         when x"B08" => Q := "111000";
         when x"B09" => Q := "111000";


-- CH=B1 
         when x"B10" => Q := "111000";
         when x"B11" => Q := "111000";
         when x"B12" => Q := "111000";
         when x"B17" => Q := "111000";
         when x"B18" => Q := "111000";
         when x"B19" => Q := "111000";


-- CH=B2 
         when x"B20" => Q := "000111";
         when x"B21" => Q := "000111";
         when x"B22" => Q := "000111";
         when x"B27" => Q := "111000";
         when x"B28" => Q := "111000";
         when x"B29" => Q := "111000";


-- CH=B3 
         when x"B30" => Q := "111111";
         when x"B31" => Q := "111111";
         when x"B32" => Q := "111111";
         when x"B37" => Q := "111000";
         when x"B38" => Q := "111000";
         when x"B39" => Q := "111000";


-- CH=B4 
         when x"B43" => Q := "111000";
         when x"B44" => Q := "111000";
         when x"B45" => Q := "111000";
         when x"B46" => Q := "111000";
         when x"B47" => Q := "111000";
         when x"B48" => Q := "111000";
         when x"B49" => Q := "111000";


-- CH=B5 
         when x"B50" => Q := "111000";
         when x"B51" => Q := "111000";
         when x"B52" => Q := "111000";
         when x"B53" => Q := "111000";
         when x"B54" => Q := "111000";
         when x"B55" => Q := "111000";
         when x"B56" => Q := "111000";
         when x"B57" => Q := "111000";
         when x"B58" => Q := "111000";
         when x"B59" => Q := "111000";


-- CH=B6 
         when x"B60" => Q := "000111";
         when x"B61" => Q := "000111";
         when x"B62" => Q := "000111";
         when x"B63" => Q := "111000";
         when x"B64" => Q := "111000";
         when x"B65" => Q := "111000";
         when x"B66" => Q := "111000";
         when x"B67" => Q := "111000";
         when x"B68" => Q := "111000";
         when x"B69" => Q := "111000";


-- CH=B7 
         when x"B70" => Q := "111111";
         when x"B71" => Q := "111111";
         when x"B72" => Q := "111111";
         when x"B73" => Q := "111000";
         when x"B74" => Q := "111000";
         when x"B75" => Q := "111000";
         when x"B76" => Q := "111000";
         when x"B77" => Q := "111000";
         when x"B78" => Q := "111000";
         when x"B79" => Q := "111000";


-- CH=B8 
         when x"B83" => Q := "000111";
         when x"B84" => Q := "000111";
         when x"B85" => Q := "000111";
         when x"B86" => Q := "000111";
         when x"B87" => Q := "111000";
         when x"B88" => Q := "111000";
         when x"B89" => Q := "111000";


-- CH=B9 
         when x"B90" => Q := "111000";
         when x"B91" => Q := "111000";
         when x"B92" => Q := "111000";
         when x"B93" => Q := "000111";
         when x"B94" => Q := "000111";
         when x"B95" => Q := "000111";
         when x"B96" => Q := "000111";
         when x"B97" => Q := "111000";
         when x"B98" => Q := "111000";
         when x"B99" => Q := "111000";


-- CH=BA 
         when x"BA0" => Q := "000111";
         when x"BA1" => Q := "000111";
         when x"BA2" => Q := "000111";
         when x"BA3" => Q := "000111";
         when x"BA4" => Q := "000111";
         when x"BA5" => Q := "000111";
         when x"BA6" => Q := "000111";
         when x"BA7" => Q := "111000";
         when x"BA8" => Q := "111000";
         when x"BA9" => Q := "111000";


-- CH=BB 
         when x"BB0" => Q := "111111";
         when x"BB1" => Q := "111111";
         when x"BB2" => Q := "111111";
         when x"BB3" => Q := "000111";
         when x"BB4" => Q := "000111";
         when x"BB5" => Q := "000111";
         when x"BB6" => Q := "000111";
         when x"BB7" => Q := "111000";
         when x"BB8" => Q := "111000";
         when x"BB9" => Q := "111000";


-- CH=BC 
         when x"BC3" => Q := "111111";
         when x"BC4" => Q := "111111";
         when x"BC5" => Q := "111111";
         when x"BC6" => Q := "111111";
         when x"BC7" => Q := "111000";
         when x"BC8" => Q := "111000";
         when x"BC9" => Q := "111000";


-- CH=BD 
         when x"BD0" => Q := "111000";
         when x"BD1" => Q := "111000";
         when x"BD2" => Q := "111000";
         when x"BD3" => Q := "111111";
         when x"BD4" => Q := "111111";
         when x"BD5" => Q := "111111";
         when x"BD6" => Q := "111111";
         when x"BD7" => Q := "111000";
         when x"BD8" => Q := "111000";
         when x"BD9" => Q := "111000";


-- CH=BE 
         when x"BE0" => Q := "000111";
         when x"BE1" => Q := "000111";
         when x"BE2" => Q := "000111";
         when x"BE3" => Q := "111111";
         when x"BE4" => Q := "111111";
         when x"BE5" => Q := "111111";
         when x"BE6" => Q := "111111";
         when x"BE7" => Q := "111000";
         when x"BE8" => Q := "111000";
         when x"BE9" => Q := "111000";


-- CH=BF 
         when x"BF0" => Q := "111111";
         when x"BF1" => Q := "111111";
         when x"BF2" => Q := "111111";
         when x"BF3" => Q := "111111";
         when x"BF4" => Q := "111111";
         when x"BF5" => Q := "111111";
         when x"BF6" => Q := "111111";
         when x"BF7" => Q := "111000";
         when x"BF8" => Q := "111000";
         when x"BF9" => Q := "111000";


-- CH=C0 
         when x"C01" => Q := "001110";
         when x"C02" => Q := "010001";
         when x"C03" => Q := "010111";
         when x"C04" => Q := "010101";
         when x"C05" => Q := "010111";
         when x"C06" => Q := "010000";
         when x"C07" => Q := "001110";


-- CH=C1 
         when x"C11" => Q := "000100";
         when x"C12" => Q := "001010";
         when x"C13" => Q := "010001";
         when x"C14" => Q := "010001";
         when x"C15" => Q := "011111";
         when x"C16" => Q := "010001";
         when x"C17" => Q := "010001";


-- CH=C2 
         when x"C21" => Q := "011110";
         when x"C22" => Q := "010001";
         when x"C23" => Q := "010001";
         when x"C24" => Q := "011110";
         when x"C25" => Q := "010001";
         when x"C26" => Q := "010001";
         when x"C27" => Q := "011110";


-- CH=C3 
         when x"C31" => Q := "001110";
         when x"C32" => Q := "010001";
         when x"C33" => Q := "010000";
         when x"C34" => Q := "010000";
         when x"C35" => Q := "010000";
         when x"C36" => Q := "010001";
         when x"C37" => Q := "001110";


-- CH=C4 
         when x"C41" => Q := "011110";
         when x"C42" => Q := "010001";
         when x"C43" => Q := "010001";
         when x"C44" => Q := "010001";
         when x"C45" => Q := "010001";
         when x"C46" => Q := "010001";
         when x"C47" => Q := "011110";


-- CH=C5 
         when x"C51" => Q := "011111";
         when x"C52" => Q := "010000";
         when x"C53" => Q := "010000";
         when x"C54" => Q := "011110";
         when x"C55" => Q := "010000";
         when x"C56" => Q := "010000";
         when x"C57" => Q := "011111";


-- CH=C6 
         when x"C61" => Q := "011111";
         when x"C62" => Q := "010000";
         when x"C63" => Q := "010000";
         when x"C64" => Q := "011110";
         when x"C65" => Q := "010000";
         when x"C66" => Q := "010000";
         when x"C67" => Q := "010000";


-- CH=C7 
         when x"C71" => Q := "001110";
         when x"C72" => Q := "010001";
         when x"C73" => Q := "010000";
         when x"C74" => Q := "010000";
         when x"C75" => Q := "010011";
         when x"C76" => Q := "010001";
         when x"C77" => Q := "001111";


-- CH=C8 
         when x"C81" => Q := "010001";
         when x"C82" => Q := "010001";
         when x"C83" => Q := "010001";
         when x"C84" => Q := "011111";
         when x"C85" => Q := "010001";
         when x"C86" => Q := "010001";
         when x"C87" => Q := "010001";


-- CH=C9 
         when x"C91" => Q := "001110";
         when x"C92" => Q := "000100";
         when x"C93" => Q := "000100";
         when x"C94" => Q := "000100";
         when x"C95" => Q := "000100";
         when x"C96" => Q := "000100";
         when x"C97" => Q := "001110";


-- CH=CA 
         when x"CA1" => Q := "000001";
         when x"CA2" => Q := "000001";
         when x"CA3" => Q := "000001";
         when x"CA4" => Q := "000001";
         when x"CA5" => Q := "000001";
         when x"CA6" => Q := "010001";
         when x"CA7" => Q := "001110";


-- CH=CB 
         when x"CB1" => Q := "010001";
         when x"CB2" => Q := "010010";
         when x"CB3" => Q := "010100";
         when x"CB4" => Q := "011000";
         when x"CB5" => Q := "010100";
         when x"CB6" => Q := "010010";
         when x"CB7" => Q := "010001";


-- CH=CC 
         when x"CC1" => Q := "010000";
         when x"CC2" => Q := "010000";
         when x"CC3" => Q := "010000";
         when x"CC4" => Q := "010000";
         when x"CC5" => Q := "010000";
         when x"CC6" => Q := "010000";
         when x"CC7" => Q := "011111";


-- CH=CD 
         when x"CD1" => Q := "010001";
         when x"CD2" => Q := "011011";
         when x"CD3" => Q := "010101";
         when x"CD4" => Q := "010101";
         when x"CD5" => Q := "010001";
         when x"CD6" => Q := "010001";
         when x"CD7" => Q := "010001";


-- CH=CE 
         when x"CE1" => Q := "010001";
         when x"CE2" => Q := "010001";
         when x"CE3" => Q := "011001";
         when x"CE4" => Q := "010101";
         when x"CE5" => Q := "010011";
         when x"CE6" => Q := "010001";
         when x"CE7" => Q := "010001";


-- CH=CF 
         when x"CF1" => Q := "001110";
         when x"CF2" => Q := "010001";
         when x"CF3" => Q := "010001";
         when x"CF4" => Q := "010001";
         when x"CF5" => Q := "010001";
         when x"CF6" => Q := "010001";
         when x"CF7" => Q := "001110";


-- CH=D0 
         when x"D01" => Q := "011110";
         when x"D02" => Q := "010001";
         when x"D03" => Q := "010001";
         when x"D04" => Q := "011110";
         when x"D05" => Q := "010000";
         when x"D06" => Q := "010000";
         when x"D07" => Q := "010000";


-- CH=D1 
         when x"D11" => Q := "001110";
         when x"D12" => Q := "010001";
         when x"D13" => Q := "010001";
         when x"D14" => Q := "010001";
         when x"D15" => Q := "010101";
         when x"D16" => Q := "010010";
         when x"D17" => Q := "001101";


-- CH=D2 
         when x"D21" => Q := "011110";
         when x"D22" => Q := "010001";
         when x"D23" => Q := "010001";
         when x"D24" => Q := "011110";
         when x"D25" => Q := "010100";
         when x"D26" => Q := "010010";
         when x"D27" => Q := "010001";


-- CH=D3 
         when x"D31" => Q := "001110";
         when x"D32" => Q := "010001";
         when x"D33" => Q := "010000";
         when x"D34" => Q := "001110";
         when x"D35" => Q := "000001";
         when x"D36" => Q := "010001";
         when x"D37" => Q := "001110";


-- CH=D4 
         when x"D41" => Q := "011111";
         when x"D42" => Q := "000100";
         when x"D43" => Q := "000100";
         when x"D44" => Q := "000100";
         when x"D45" => Q := "000100";
         when x"D46" => Q := "000100";
         when x"D47" => Q := "000100";


-- CH=D5 
         when x"D51" => Q := "010001";
         when x"D52" => Q := "010001";
         when x"D53" => Q := "010001";
         when x"D54" => Q := "010001";
         when x"D55" => Q := "010001";
         when x"D56" => Q := "010001";
         when x"D57" => Q := "001110";


-- CH=D6 
         when x"D61" => Q := "010001";
         when x"D62" => Q := "010001";
         when x"D63" => Q := "010001";
         when x"D64" => Q := "001010";
         when x"D65" => Q := "001010";
         when x"D66" => Q := "000100";
         when x"D67" => Q := "000100";


-- CH=D7 
         when x"D71" => Q := "010001";
         when x"D72" => Q := "010001";
         when x"D73" => Q := "010001";
         when x"D74" => Q := "010101";
         when x"D75" => Q := "010101";
         when x"D76" => Q := "010101";
         when x"D77" => Q := "001010";


-- CH=D8 
         when x"D81" => Q := "010001";
         when x"D82" => Q := "010001";
         when x"D83" => Q := "001010";
         when x"D84" => Q := "000100";
         when x"D85" => Q := "001010";
         when x"D86" => Q := "010001";
         when x"D87" => Q := "010001";


-- CH=D9 
         when x"D91" => Q := "010001";
         when x"D92" => Q := "010001";
         when x"D93" => Q := "001010";
         when x"D94" => Q := "000100";
         when x"D95" => Q := "000100";
         when x"D96" => Q := "000100";
         when x"D97" => Q := "000100";


-- CH=DA 
         when x"DA1" => Q := "011111";
         when x"DA2" => Q := "000001";
         when x"DA3" => Q := "000010";
         when x"DA4" => Q := "000100";
         when x"DA5" => Q := "001000";
         when x"DA6" => Q := "010000";
         when x"DA7" => Q := "011111";


-- CH=DB 
         when x"DB2" => Q := "000100";
         when x"DB3" => Q := "001000";
         when x"DB4" => Q := "011111";
         when x"DB5" => Q := "001000";
         when x"DB6" => Q := "000100";


-- CH=DC 
         when x"DC1" => Q := "010000";
         when x"DC2" => Q := "010000";
         when x"DC3" => Q := "010000";
         when x"DC4" => Q := "010000";
         when x"DC5" => Q := "010110";
         when x"DC6" => Q := "000001";
         when x"DC7" => Q := "000010";
         when x"DC8" => Q := "000100";
         when x"DC9" => Q := "000111";


-- CH=DD 
         when x"DD2" => Q := "000100";
         when x"DD3" => Q := "000010";
         when x"DD4" => Q := "011111";
         when x"DD5" => Q := "000010";
         when x"DD6" => Q := "000100";


-- CH=DE 
         when x"DE2" => Q := "000100";
         when x"DE3" => Q := "001110";
         when x"DE4" => Q := "010101";
         when x"DE5" => Q := "000100";
         when x"DE6" => Q := "000100";


-- CH=DF 
         when x"DF1" => Q := "001010";
         when x"DF2" => Q := "001010";
         when x"DF3" => Q := "011111";
         when x"DF4" => Q := "001010";
         when x"DF5" => Q := "011111";
         when x"DF6" => Q := "001010";
         when x"DF7" => Q := "001010";


-- CH=E0 
         when x"E07" => Q := "000111";
         when x"E08" => Q := "000111";
         when x"E09" => Q := "000111";


-- CH=E1 
         when x"E10" => Q := "111000";
         when x"E11" => Q := "111000";
         when x"E12" => Q := "111000";
         when x"E17" => Q := "000111";
         when x"E18" => Q := "000111";
         when x"E19" => Q := "000111";


-- CH=E2 
         when x"E20" => Q := "000111";
         when x"E21" => Q := "000111";
         when x"E22" => Q := "000111";
         when x"E27" => Q := "000111";
         when x"E28" => Q := "000111";
         when x"E29" => Q := "000111";


-- CH=E3 
         when x"E30" => Q := "111111";
         when x"E31" => Q := "111111";
         when x"E32" => Q := "111111";
         when x"E37" => Q := "000111";
         when x"E38" => Q := "000111";
         when x"E39" => Q := "000111";


-- CH=E4 
         when x"E43" => Q := "111000";
         when x"E44" => Q := "111000";
         when x"E45" => Q := "111000";
         when x"E46" => Q := "111000";
         when x"E47" => Q := "000111";
         when x"E48" => Q := "000111";
         when x"E49" => Q := "000111";


-- CH=E5 
         when x"E50" => Q := "111000";
         when x"E51" => Q := "111000";
         when x"E52" => Q := "111000";
         when x"E53" => Q := "111000";
         when x"E54" => Q := "111000";
         when x"E55" => Q := "111000";
         when x"E56" => Q := "111000";
         when x"E57" => Q := "000111";
         when x"E58" => Q := "000111";
         when x"E59" => Q := "000111";


-- CH=E6 
         when x"E60" => Q := "000111";
         when x"E61" => Q := "000111";
         when x"E62" => Q := "000111";
         when x"E63" => Q := "111000";
         when x"E64" => Q := "111000";
         when x"E65" => Q := "111000";
         when x"E66" => Q := "111000";
         when x"E67" => Q := "000111";
         when x"E68" => Q := "000111";
         when x"E69" => Q := "000111";


-- CH=E7 
         when x"E70" => Q := "111111";
         when x"E71" => Q := "111111";
         when x"E72" => Q := "111111";
         when x"E73" => Q := "111000";
         when x"E74" => Q := "111000";
         when x"E75" => Q := "111000";
         when x"E76" => Q := "111000";
         when x"E77" => Q := "000111";
         when x"E78" => Q := "000111";
         when x"E79" => Q := "000111";


-- CH=E8 
         when x"E83" => Q := "000111";
         when x"E84" => Q := "000111";
         when x"E85" => Q := "000111";
         when x"E86" => Q := "000111";
         when x"E87" => Q := "000111";
         when x"E88" => Q := "000111";
         when x"E89" => Q := "000111";


-- CH=E9 
         when x"E90" => Q := "111000";
         when x"E91" => Q := "111000";
         when x"E92" => Q := "111000";
         when x"E93" => Q := "000111";
         when x"E94" => Q := "000111";
         when x"E95" => Q := "000111";
         when x"E96" => Q := "000111";
         when x"E97" => Q := "000111";
         when x"E98" => Q := "000111";
         when x"E99" => Q := "000111";


-- CH=EA 
         when x"EA0" => Q := "000111";
         when x"EA1" => Q := "000111";
         when x"EA2" => Q := "000111";
         when x"EA3" => Q := "000111";
         when x"EA4" => Q := "000111";
         when x"EA5" => Q := "000111";
         when x"EA6" => Q := "000111";
         when x"EA7" => Q := "000111";
         when x"EA8" => Q := "000111";
         when x"EA9" => Q := "000111";


-- CH=EB 
         when x"EB0" => Q := "111111";
         when x"EB1" => Q := "111111";
         when x"EB2" => Q := "111111";
         when x"EB3" => Q := "000111";
         when x"EB4" => Q := "000111";
         when x"EB5" => Q := "000111";
         when x"EB6" => Q := "000111";
         when x"EB7" => Q := "000111";
         when x"EB8" => Q := "000111";
         when x"EB9" => Q := "000111";


-- CH=EC 
         when x"EC3" => Q := "111111";
         when x"EC4" => Q := "111111";
         when x"EC5" => Q := "111111";
         when x"EC6" => Q := "111111";
         when x"EC7" => Q := "000111";
         when x"EC8" => Q := "000111";
         when x"EC9" => Q := "000111";


-- CH=ED 
         when x"ED0" => Q := "111000";
         when x"ED1" => Q := "111000";
         when x"ED2" => Q := "111000";
         when x"ED3" => Q := "111111";
         when x"ED4" => Q := "111111";
         when x"ED5" => Q := "111111";
         when x"ED6" => Q := "111111";
         when x"ED7" => Q := "000111";
         when x"ED8" => Q := "000111";
         when x"ED9" => Q := "000111";


-- CH=EE 
         when x"EE0" => Q := "000111";
         when x"EE1" => Q := "000111";
         when x"EE2" => Q := "000111";
         when x"EE3" => Q := "111111";
         when x"EE4" => Q := "111111";
         when x"EE5" => Q := "111111";
         when x"EE6" => Q := "111111";
         when x"EE7" => Q := "000111";
         when x"EE8" => Q := "000111";
         when x"EE9" => Q := "000111";


-- CH=EF 
         when x"EF0" => Q := "111111";
         when x"EF1" => Q := "111111";
         when x"EF2" => Q := "111111";
         when x"EF3" => Q := "111111";
         when x"EF4" => Q := "111111";
         when x"EF5" => Q := "111111";
         when x"EF6" => Q := "111111";
         when x"EF7" => Q := "000111";
         when x"EF8" => Q := "000111";
         when x"EF9" => Q := "000111";


-- CH=F0 
         when x"F07" => Q := "111111";
         when x"F08" => Q := "111111";
         when x"F09" => Q := "111111";


-- CH=F1 
         when x"F10" => Q := "111000";
         when x"F11" => Q := "111000";
         when x"F12" => Q := "111000";
         when x"F17" => Q := "111111";
         when x"F18" => Q := "111111";
         when x"F19" => Q := "111111";


-- CH=F2 
         when x"F20" => Q := "000111";
         when x"F21" => Q := "000111";
         when x"F22" => Q := "000111";
         when x"F27" => Q := "111111";
         when x"F28" => Q := "111111";
         when x"F29" => Q := "111111";


-- CH=F3 
         when x"F30" => Q := "111111";
         when x"F31" => Q := "111111";
         when x"F32" => Q := "111111";
         when x"F37" => Q := "111111";
         when x"F38" => Q := "111111";
         when x"F39" => Q := "111111";


-- CH=F4 
         when x"F43" => Q := "111000";
         when x"F44" => Q := "111000";
         when x"F45" => Q := "111000";
         when x"F46" => Q := "111000";
         when x"F47" => Q := "111111";
         when x"F48" => Q := "111111";
         when x"F49" => Q := "111111";


-- CH=F5 
         when x"F50" => Q := "111000";
         when x"F51" => Q := "111000";
         when x"F52" => Q := "111000";
         when x"F53" => Q := "111000";
         when x"F54" => Q := "111000";
         when x"F55" => Q := "111000";
         when x"F56" => Q := "111000";
         when x"F57" => Q := "111111";
         when x"F58" => Q := "111111";
         when x"F59" => Q := "111111";


-- CH=F6 
         when x"F60" => Q := "000111";
         when x"F61" => Q := "000111";
         when x"F62" => Q := "000111";
         when x"F63" => Q := "111000";
         when x"F64" => Q := "111000";
         when x"F65" => Q := "111000";
         when x"F66" => Q := "111000";
         when x"F67" => Q := "111111";
         when x"F68" => Q := "111111";
         when x"F69" => Q := "111111";


-- CH=F7 
         when x"F70" => Q := "111111";
         when x"F71" => Q := "111111";
         when x"F72" => Q := "111111";
         when x"F73" => Q := "111000";
         when x"F74" => Q := "111000";
         when x"F75" => Q := "111000";
         when x"F76" => Q := "111000";
         when x"F77" => Q := "111111";
         when x"F78" => Q := "111111";
         when x"F79" => Q := "111111";


-- CH=F8 
         when x"F83" => Q := "000111";
         when x"F84" => Q := "000111";
         when x"F85" => Q := "000111";
         when x"F86" => Q := "000111";
         when x"F87" => Q := "111111";
         when x"F88" => Q := "111111";
         when x"F89" => Q := "111111";


-- CH=F9 
         when x"F90" => Q := "111000";
         when x"F91" => Q := "111000";
         when x"F92" => Q := "111000";
         when x"F93" => Q := "000111";
         when x"F94" => Q := "000111";
         when x"F95" => Q := "000111";
         when x"F96" => Q := "000111";
         when x"F97" => Q := "111111";
         when x"F98" => Q := "111111";
         when x"F99" => Q := "111111";


-- CH=FA 
         when x"FA0" => Q := "000111";
         when x"FA1" => Q := "000111";
         when x"FA2" => Q := "000111";
         when x"FA3" => Q := "000111";
         when x"FA4" => Q := "000111";
         when x"FA5" => Q := "000111";
         when x"FA6" => Q := "000111";
         when x"FA7" => Q := "111111";
         when x"FA8" => Q := "111111";
         when x"FA9" => Q := "111111";


-- CH=FB 
         when x"FB0" => Q := "111111";
         when x"FB1" => Q := "111111";
         when x"FB2" => Q := "111111";
         when x"FB3" => Q := "000111";
         when x"FB4" => Q := "000111";
         when x"FB5" => Q := "000111";
         when x"FB6" => Q := "000111";
         when x"FB7" => Q := "111111";
         when x"FB8" => Q := "111111";
         when x"FB9" => Q := "111111";


-- CH=FC 
         when x"FC3" => Q := "111111";
         when x"FC4" => Q := "111111";
         when x"FC5" => Q := "111111";
         when x"FC6" => Q := "111111";
         when x"FC7" => Q := "111111";
         when x"FC8" => Q := "111111";
         when x"FC9" => Q := "111111";


-- CH=FD 
         when x"FD0" => Q := "111000";
         when x"FD1" => Q := "111000";
         when x"FD2" => Q := "111000";
         when x"FD3" => Q := "111111";
         when x"FD4" => Q := "111111";
         when x"FD5" => Q := "111111";
         when x"FD6" => Q := "111111";
         when x"FD7" => Q := "111111";
         when x"FD8" => Q := "111111";
         when x"FD9" => Q := "111111";


-- CH=FE 
         when x"FE0" => Q := "000111";
         when x"FE1" => Q := "000111";
         when x"FE2" => Q := "000111";
         when x"FE3" => Q := "111111";
         when x"FE4" => Q := "111111";
         when x"FE5" => Q := "111111";
         when x"FE6" => Q := "111111";
         when x"FE7" => Q := "111111";
         when x"FE8" => Q := "111111";
         when x"FE9" => Q := "111111";


-- CH=FF 
         when x"FF0" => Q := "111111";
         when x"FF1" => Q := "111111";
         when x"FF2" => Q := "111111";
         when x"FF3" => Q := "111111";
         when x"FF4" => Q := "111111";
         when x"FF5" => Q := "111111";
         when x"FF6" => Q := "111111";
         when x"FF7" => Q := "111111";
         when x"FF8" => Q := "111111";
         when x"FF9" => Q := "111111";

	   	when others => Q := (others => '0');

	   end case;

	   TOP := A(11) and A(9);

	   if r_switch = '0' then
	   	QA <= TOP & "0" & Q;
	   else
	   	QB <= TOP & "0" & Q;
	   end if;

		r_switch <= not r_switch;
	end if;

end process;

end RTL;